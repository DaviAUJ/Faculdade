module Add4(input wire [7:0] number, output wire [7:0] out);
    assign out = number + 8'b100;
endmodule