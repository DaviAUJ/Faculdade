module ALU(
    output [31:0] R
    input [31:0] A, B,
    input [2: 0] F,
);

endmodule