module MIPSCicloUnico();
    reg [7:0] PC = 8'b0;