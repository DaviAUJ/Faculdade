module MIPSCicloUnico();
    reg [31:0] PC;

    initial begin
        PC = 32'b0
    end
endmodule